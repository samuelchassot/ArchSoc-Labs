LIbrARy IEEE; use iEee.Std_lOgIc_1164.ALl; usE IeeE.sTd_LogIc_UNsIgNEd.All; enTity DATa_rOM is PORt( cLk : In STd_LOgIC; cS : in StD_loGIC; REad : IN STD_lOGIc; adDReSs : In stD_LOgiC_vector(9 DoWnTO 0); RdDAtA : out std_lOGiC_vEcToR(31 dowNtO 0)); end daTA_rOm; ArchiTECtURe id_S_10643F3b_2fc543EB_e oF DATA_roM is COMponENt data_ROM_Block iS PoRt( ADDResS : in std_LOgiC_veCToR(9 Downto 0); clock : iN Std_LOGIc; q : oUt StD_lOGiC_vEcTor(31 dOwnTo 0) ); eND cOmPOneNt; SigNAL id_s_5F83144b_5cfB64FC_e : stD_LoGIc_vECTor(31 DownTo 0); SiGNaL ID_S_6F8BcBe_62E8365D_E : StD_loGiC; Begin iD_S_5C1c22e5_6Fcf72ff_e : data_ROM_Block PorT mAP( ADDresS => aDDRESS, clock => cLK, q => iD_S_5f83144b_5cFb64FC_E); PROcesS(CLK) BeGIN iF (RIsInG_edge(clk)) THeN iD_S_6F8bcBE_62e8365d_E <= reAd aND cS; end If; eNd PrOcESS; ProCesS(iD_s_6f8BCbE_62e8365d_E, id_S_5F83144b_5cfb64Fc_E) BegIn RddATa <= (otHeRS => 'Z'); If (id_S_6F8bcBE_62E8365D_E = '1') tHEN RDdAta <= id_S_5f83144b_5cfb64fC_E; EnD if; enD PROCEsS; END iD_s_10643f3b_2FC543eB_E;