LIBRARY IeEE; use IeEe.stD_LOgIc_1164.ALl; usE ieEE.StD_LOgIC_uNSIgNED.aLL; ENtity iNStrUctiOn_RoM iS POrt( ClK : In sTD_LOgic; cS : iN stD_loGIC; rEaD : iN STd_logiC; addREss : In StD_LogIC_VeCTOr(9 DOwNtO 0); rddaTa : out sTd_LoGic_VECToR(31 DOwNTo 0)); End iNStRUCtion_ROm; aRchiTEcTUrE id_S_10643F3b_2FC543EB_e OF InsTRUctIOn_rOM iS cOMPONENT instruction_ROM_Block is POrt( aDDrEss : in StD_LOgIC_VectOr(9 dowNTo 0); clock : iN StD_LogIC; q : OuT std_lOGic_vEcToR(31 dOwnTo 0) ); END coMponent; sIgnAl ID_S_5F83144B_5cFb64FC_e : STd_LOgIC_VECTOR(31 dOwnto 0); siGNAl iD_s_6F8bcbe_62e8365d_e : STD_lOgIc; BeGIn iD_S_36FDD56D_59c20fa9_E : instruction_ROM_Block pORt MAP( aDdreSS => aDDrEss, clock => Clk, q => iD_s_5f83144b_5cFB64FC_e); PRoceSS(clK) Begin if (rISiNG_EdGe(cLK)) THeN id_s_6f8Bcbe_62E8365D_e <= READ aND cs; EnD IF; ENd pRocESs; PROcESS(id_S_6F8bCBe_62E8365d_E, iD_S_5F83144b_5Cfb64Fc_e) begIn rdDatA <= (otHERs => 'Z'); IF (iD_s_6f8bcbe_62E8365d_E = '1') theN RddATa <= iD_s_5f83144b_5CFB64fc_e; END If; End prOcess; end ID_s_10643F3B_2fc543eB_e;